----------------------------------------------------------------------------------
-- MOBY-DIC Project
-- www.mobydic-project.eu
--
-- Copyright:
-- (C) 2011 Tomaso Poggi, Spain, tpoggi@essbilbao.org
-- (C) 2011 Alberto Oliveri, University of Genoa, Italy, alberto.oliveri@unige.it
--
-- Legal note:
-- This program is free software; you can redistribute it and/or
-- modify it under the terms of the GNU General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License, or (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- General Public License for more details.
-- 
-- You should have received a copy of the GNU General Public
-- License along with this library; if not, write to the 
-- Free Software Foundation, Inc., 
-- 59 Temple Place, Suite 330, 
-- Boston, MA  02111-1307  USA
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.pwasFunctionPackage.all;

entity Memory is
	Port ( clk : in std_logic;
	     start : in std_logic;
	     reset : in std_logic;
	      addr : in addr_matrix_pwas;
	       res : out mem_matrix_pwas;
	      done : out std_logic);
end Memory;

-- Architecture declaration

architecture Behavioral of Memory is
		
--- BEGIN MATLABGEN ---

	type ROM_type is array (0 to 5119) of signed(N_BIT_COEFF_PWAS-1 downto 0);

	constant ROM_0 : ROM_type:=(
	"001000111110", "111011110010", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111110110", "100010110011", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "000111100111", "011010001010", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"000111011010", "000111011010", "001010100100", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001001000011", "001010001010", "001010000111", "001010000100", "001010001000", "001100110111", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000011110001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100010000", "111100000010", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111110101", "100011101100", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"000111011010", "011010001010", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011100", "010010010001", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111101001", "000111011010", "000111011010", "001000000111", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000010010011", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001001001110", "111101010011", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111101100", 
	"100011001111", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111100000", "011010010000", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "000111011010", "000111011010", "001011010010", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001000110011", "001001101010", "001001100100", "001001100100", 
	"001001100101", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000011001001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001011111111", "111111111111", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "100011101100", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "000111011010", "011010010000", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", 
	"010010110001", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "000111011010", "001100101101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000001001001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001001001101", "111101010101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111101100", "100011001111", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111100000", "011010010000", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "001011010001", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001000110100", "001001101101", 
	"001001100111", "001001101000", "001001100111", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000011001001", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001011111110", "111111111111", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "100011101100", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "011010010000", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"000111011010", "000111011010", "010010110010", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "000111011010", "001100110111", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000001001001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001001001101", "111101010101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111101100", "100011001111", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"000111100000", "011010010000", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "001011010001", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001000110100", "001001101101", "001001100111", "001001100111", "001001100110", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000011001001", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001011111110", "111111111111", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"100011101100", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "011010010000", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "000111011010", "000111011010", "010010110010", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", 
	"000111011010", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000001001001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001001001101", "111101010101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111101100", "100011001111", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "000111100000", "011010010000", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", 
	"001011010001", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001000110100", "001001101101", "001001100111", "001001101000", "001001100111", "001100110111", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000011001001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001011111110", "111111111111", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "100011101100", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "011010010000", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "010010110010", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"000111011010", "000111011010", "000111011010", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000001001001", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001001001101", "111101010101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111101100", "100011001111", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "000111100000", "011010010000", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"000111011010", "000111011010", "001011010001", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001000110100", "001001101101", "001001100111", "001001101000", "001001100111", "001100110111", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000011001001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001011111110", "111111111111", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "100011101100", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"000111011010", "011010010000", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "010010110010", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "000111011010", "000111011010", "000111011010", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000001001001", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001001001101", "111101010101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111101100", 
	"100011001111", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111100000", "011010010000", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "000111011010", "000111011010", "001011010001", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001000110100", "001001101101", "001001100111", "001001101000", 
	"001001100111", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000011001001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001011111110", "111111111111", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "100011101100", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "000111011010", "011010010000", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", 
	"010010110010", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "000111011010", "001100110111", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000001001001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001001001110", "111101010001", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111101100", "100011001111", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111100000", "011010010000", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "001011010000", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001000110011", "001001101011", 
	"001001100110", "001001100111", "001001100110", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000011001001", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001011111110", "111111111111", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "100011101100", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "011010010000", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"000111011010", "000111011010", "010010110010", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "000111011010", "001100110111", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000001001001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001000111101", "111100110110", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111101100", "100011001111", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"000111100000", "011010010000", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "001011101110", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001001000011", "001001111010", "001001110100", "001001110100", "001001101011", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000011001001", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001100000000", "111111111111", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"100011101100", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "011010010000", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "000111011010", "000111011010", "010010110010", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", 
	"000111011010", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000001001001", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100011100", "111100110110", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111101111", "100011101011", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "000111011010", "011010010000", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", 
	"010010010010", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111101110", "000111100010", "000111100010", "001000000110", "001100110111", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000010010011", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000101100101", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001100010001", "111111111111", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000111011010", "000111011010", "100011101100", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "011010010000", 
	"000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000111011010", "000111011010", "000111011010", "000111011010", "010101010111", "000101100101", "000101100101", "000101100101", 
	"000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000111011010", "000111011010", 
	"000111011010", "000111011010", "000111011010", "001100110111", "000101100101", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "001100100010", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "000101100101", "000101100101", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000101100101", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000101100101", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000101100101", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", 
	"001100110111", "001100110111", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000101100101", "000101100101", 
	"001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "001100110111", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", 
	"000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000", "000000000000");

begin

	proc_mem: process(clk,reset)
	begin
		if reset = '0' then
			for i in 0 to N_FUN_PWAS-1 loop
				for j in 0 to N_DIM_PWAS loop
					res(i)(j) <= (others => '0');
				end loop;
			end loop;
		elsif rising_edge(clk) and start = '1' then
			for j in 0 to N_DIM_PWAS loop
				res(0)(j) <= '0'&ROM_0(to_integer(addr(j)));
			end loop;
		end if;
	end process;
--- END MATLABGEN ---
	
	done <= '0' when reset = '0' else
	        start when rising_edge(clk);
	

end Behavioral;
