--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package pwagFunctionPackage is

	-- Declare constants
	
--- BEGIN MATLABGEN ---
--- END MATLABGEN ---

end pwagFunctionPackage;
