----------------------------------------------------------------------------------
-- MOBY-DIC Project
-- www.mobydic-project.eu
--
-- Copyright:
-- (C) 2011 Tomaso Poggi, Spain, tpoggi@essbilbao.org
-- (C) 2011 Alberto Oliveri, University of Genoa, Italy, alberto.oliveri@unige.it
--
-- Legal note:
-- This program is free software; you can redistribute it and/or
-- modify it under the terms of the GNU General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License, or (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- General Public License for more details.
-- 
-- You should have received a copy of the GNU General Public
-- License along with this library; if not, write to the 
-- Free Software Foundation, Inc., 
-- 59 Temple Place, Suite 330, 
-- Boston, MA  02111-1307  USA
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.pwasFunctionPackage.all;

entity Memory is
	Port ( clk : in std_logic;
	     start : in std_logic;
	     reset : in std_logic;
	      addr : in addr_matrix_pwas;
	       res : out mem_matrix_pwas;
	      done : out std_logic);
end Memory;

-- Architecture declaration

architecture Behavioral of Memory is
		
--- BEGIN MATLABGEN ---

	type ROM_type is array (0 to 63) of signed(N_BIT_COEFF_PWAS-1 downto 0);

	constant ROM_0 : ROM_type:=(
	"011111111111", "011111111111", "011111111111", "011111111111", "011111111101", "011111111101", "011111111101", "011111111100", "011111111111", "011111111111", 
	"011111111111", "011111111101", "011111111110", "011111111110", "011111111110", "011111111110", "011111111111", "011111111111", "011111111101", "011111111111", 
	"011111111111", "011111111111", "011111111111", "011111111111", "011111111111", "011111111111", "011111111111", "011111111111", "001110100111", "111101000100", 
	"101100001010", "100000000000", "011111111111", "001101001000", "111011010000", "101000010010", "100000000000", "100000000000", "100000000000", "100000000000", 
	"100010011100", "100000000000", "100000000000", "100000000000", "100000000000", "100000000001", "100000000001", "100000000000", "100000000000", "100000000000", 
	"100000000001", "100000000001", "100000000001", "100000000001", "100000000000", "100000000000", "100000000011", "100000000010", "100000000010", "100000000010", 
	"100000000010", "100000000000", "100000000000", "100000000000");

begin

	proc_mem: process(clk,reset)
	begin
		if reset = '0' then
			for i in 0 to N_FUN_PWAS-1 loop
				for j in 0 to N_DIM_PWAS loop
					res(i)(j) <= (others => '0');
				end loop;
			end loop;
		elsif rising_edge(clk) and start = '1' then
			for j in 0 to N_DIM_PWAS loop
				res(0)(j) <= ROM_0(to_integer(addr(j)));
			end loop;
		end if;
	end process;
--- END MATLABGEN ---
	
	done <= '0' when reset = '0' else
	        start when rising_edge(clk);
	

end Behavioral;
